`default_nettype none

module system_top_level ();

endmodule
