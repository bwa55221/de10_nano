`timescale 1ns/1ps

module tb_st_sink ();



endmodule